module BUFG (
	input I,
	output O
);
	assign O = I;

endmodule
