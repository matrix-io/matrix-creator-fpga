module uart_fsm (
  input clk,    // Clock
  input resetn,  // Asynchronous reset active low
  
);





endmodule