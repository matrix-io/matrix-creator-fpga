/*
 * Copyright 2016 <Admobilize>
 * MATRIX Labs  [http://creator.matrix.one]
 * This file is part of MATRIX Creator HDL for Spartan 6
 *
 * MATRIX Creator HDL is like free software: you can redistribute 
 * it and/or modify it under the terms of the GNU General Public License 
 * as published by the Free Software Foundation, either version 3 of the 
 * License, or (at your option) any later version.

 * This program is distributed in the hope that it will be useful, but 
 * WITHOUT ANY WARRANTY; without even the implied warranty of 
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU 
 * General Public License for more details.

 * You should have received a copy of the GNU General Public License along
 * with this program.  If not, see <http://www.gnu.org/licenses/>.
 */

module core_clk#(
      parameter PRESCALER = 16
)(
      input clk,
      input rst,

      output reg [PRESCALER-1:0] core_clk);

initial begin
core_clk = 0;
end

always @(posedge clk or posedge rst ) begin
  if (rst) 
    core_clk <= 0;
  else 
    core_clk <= core_clk + 1;
end

endmodule
